library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

Library xpm;
use xpm.vcomponents.all;  -- contains clock domain crossing macros

-- This entity is a simple wrapper for the STUDENT_AREA entity,
--   providing I/Os to the board's LEDs, switches, and 
--   pushbuttons, debounced and clock-synchronised when needed.
-- It also includes a SPI_MASTER component that interfaces with
--  an external SRAM, plus the synchronisation logic required
--  to instantiate a handshaking protocol between the SPI_MASTER
--  and the STUDENT_AREA entities. 

entity TOP_LEVEL is
  Generic (disp_delay : natural := 62500000);
  Port ( 
    GCLK : in  STD_LOGIC; -- 125MHz clock
    --   BTN(0) - is wired to global reset			  
    BTN : in  STD_LOGIC_VECTOR (3 downto 0);
    -- Board switches
    SW : in  STD_LOGIC_VECTOR (1 downto 0);
    -- Board LEDs
    LED : out  STD_LOGIC_VECTOR (3 downto 0);
    -- Signals for SPI interface to SRAM
    --   Clock generated by SPI master
    SPI_SCK: out STD_LOGIC;
    --   Chip select (inverted)
    SPI_CS_INV: out STD_LOGIC;
    --   Hold signal (inverted) - not used, set to high
    SPI_HOLD_INV: out STD_LOGIC;
    --   Master-Out Slave-In serial data line
    SPI_MOSI: out STD_LOGIC;
    --   Master-In Slave-Out serial data line
    SPI_MISO: in STD_LOGIC
 );
end TOP_LEVEL;

architecture Behavioral of TOP_LEVEL is

-- Internal clock signals
signal CLK_26MHZ, CLK_125MHZ : STD_LOGIC;

-- Debounced button inputs
signal btn_db_26MHz, btn_db_125MHz : STD_LOGIC_VECTOR (3 downto 0); 

-- LED output - internal for observation
signal LD_INT : STD_LOGIC_VECTOR (3 downto 0); 

-- SWITCHES encoding (expanding from 2 to 8 bits)
signal SW_INT : STD_LOGIC_VECTOR (7 downto 0); 

-- SPI data and control signals - internal for observation
signal spi_sck_int, spi_cs_inv_int, spi_hold_inv_int, 
       spi_mosi_int, spi_miso_int : STD_LOGIC;

-- Signals to enable the SPI interface
signal en_spi, en_spi_sync: STD_LOGIC;

-- Handshaking signals for SPI write operations
signal spi_wr_ack, spi_wr_ack_sync :  STD_LOGIC;
signal spi_wr_req, spi_wr_req_sync : STD_LOGIC;

-- Handshaking signals for SPI read operations
signal spi_rd_ack, spi_rd_ack_sync :  STD_LOGIC;
signal spi_rd_req, spi_rd_req_sync : STD_LOGIC;

-- Data to/from the SPI interface
signal pdata_to_spi, pdata_from_spi : STD_LOGIC_VECTOR(7 downto 0);

-- Attributes to enable observation of internal signals
--   through the ChipScope ILA
-- UNCOMMENT TO USE ILA
attribute keep : string;
attribute keep of btn_db_26MHz : signal is "true";
attribute keep of btn_db_125MHz : signal is "true";
attribute keep of LD_INT : signal is "true";
attribute keep of spi_sck_int : signal is "true";
attribute keep of spi_cs_inv_int : signal is "true";
attribute keep of spi_hold_inv_int : signal is "true";
attribute keep of spi_mosi_int : signal is "true";
attribute keep of spi_miso_int : signal is "true";
attribute keep of en_spi : signal is "true";
attribute keep of en_spi_sync : signal is "true";
attribute keep of spi_wr_ack : signal is "true";
attribute keep of spi_wr_ack_sync : signal is "true";
attribute keep of spi_wr_req : signal is "true";
attribute keep of spi_wr_req_sync : signal is "true";
attribute keep of spi_rd_ack : signal is "true";
attribute keep of spi_rd_ack_sync : signal is "true";
attribute keep of spi_rd_req : signal is "true";
attribute keep of spi_rd_req_sync : signal is "true";
attribute keep of pdata_to_spi : signal is "true";
attribute keep of pdata_from_spi : signal is "true";


begin

-- Word to be stored in memory as a function of the
--  switch values
with SW select 
    SW_INT <= "00100100"  when "00",
              "01011010"  when "01",
              "10100101"  when "10",
              "11110001"  when "11",
              (others => 'U')    when others;
                  
-- Clock management unit: generates two clocks:
--   - 125MHz for the control logic
--   - 26MHZ for the SPI master unit
Clock_generator : entity work.CLK_GEN
port map
	(-- Clock in ports
	CLK_IN1 => GCLK,
	-- Clock out ports
	CLK_OUT1 => CLK_125MHZ,
	CLK_OUT2 => CLK_26MHZ
);

-- For the follwowing units, the input signals go through
--   two debouncers/synchronisers in series: first they 
--   are synchronised to the (slower) SPI clock, then to
--   the (faster) output clock. This ensures that each will
--   have a one-pulse duration for either clock domain and
--   that the delay between pulses is constant.

-- Debouncers and synchronisers for the (active high) user buttons. 
-- The outputs will be active-high and synchronous to the target clocks.
-- NOTE: technically they are not all needed but are left in for future
--  development (unused elements will be removed by synthesis)
debouncers: for i in 0 to 3 generate
	button_debouncer_26MHZ : entity work.Debouncer 
	PORT MAP(
		CLK => CLK_26MHZ,
		Sig => BTN(i),
		Deb_Sig => btn_db_26MHZ(i) 
	);
	button_debouncer_125_MHZ : entity work.Debouncer 
	PORT MAP(
		CLK => CLK_125MHZ,
		Sig => btn_db_26MHZ(i),
		Deb_Sig => btn_db_125MHZ(i) 
	);
end generate;

-- This entity will contain the work to be carried out for each task. 
-- Note that some I/Os might not be needed (implementation dependent)	
STUDENT_AREA_component: entity work.STUDENT_AREA 
GENERIC MAP (disp_delay => disp_delay)
PORT MAP(
    CLK => CLK_125MHZ,
    RST => btn_db_125MHZ(0), -- Note: PB(0) reserced for reset (BTND) 
    USER_PB => btn_db_125MHZ,
    SWITCHES => SW_INT,
    LEDS => LD_INT,
    DATA_FROM_SPI => pdata_from_spi,
    DATA_TO_SPI => pdata_to_spi,
    EN_SPI => en_spi,
    SPI_WR_REQ => spi_wr_req,
    SPI_WR_ACK => spi_wr_ack_sync,
    SPI_RD_REQ => spi_rd_req,
    SPI_RD_ACK => spi_rd_ack_sync,
    SRAM_ADDRESS => x"01AA05"    -- hard-wired read/write address
);

-- Cross-domain synchronisers for the handshaking and control signals
-- Note: The input data must be sampled two or more times by the 
--  destination clock

-- Enable signal for the SPI interface. Should be asserted
--  at the start of the transfer and kept high until the
--  acknowledgment for the last byte to be read is received
Sync_en_spi: xpm_cdc_single
GENERIC MAP (
  DEST_SYNC_FF => 2,   -- integer; range: 2-10
  SIM_ASSERT_CHK => 0, -- integer; 0=disable simulation messages, 
                       --          1=enable simulation messages
  SRC_INPUT_REG => 0   -- integer; 0=do not register input, 
                       --          1=register input
)
PORT MAP (
  src_clk => CLK_125MHZ,    -- used only when SRC_INPUT_REG = 1
  src_in => en_spi, 
  dest_clk => CLK_26MHZ,
  dest_out => en_spi_sync
);

-- SPI write requests generated by the output control logic
Sync_spi_wr_req: xpm_cdc_single
GENERIC MAP (
  DEST_SYNC_FF => 2,   -- integer; range: 2-10
  SIM_ASSERT_CHK => 0, -- integer; 0=disable simulation messages, 
                       --          1=enable simulation messages
  SRC_INPUT_REG => 0   -- integer; 0=do not register input, 
                       --          1=register input
)
PORT MAP (
  src_clk => CLK_125MHZ,    -- used only when SRC_INPUT_REG = 1
  src_in => spi_wr_req, 
  dest_clk => CLK_26MHZ,
  dest_out => spi_wr_req_sync
);

-- Acknowledgment of completion of a SPI write request
Sync_spi_wr_ack: xpm_cdc_single
GENERIC MAP (
  DEST_SYNC_FF => 2,   -- integer; range: 2-10
  SIM_ASSERT_CHK => 0, -- integer; 0=disable simulation messages, 
                       --          1=enable simulation messages
  SRC_INPUT_REG => 0   -- integer; 0=do not register input, 
                       --          1=register input
)
PORT MAP (
  src_clk => CLK_26MHZ,    -- used only when SRC_INPUT_REG = 1
  src_in => spi_wr_ack, 
  dest_clk => CLK_125MHZ,
  dest_out => spi_wr_ack_sync
);
			 
-- SPI read requests generated by the output control logic
Sync_spi_rd_req: xpm_cdc_single
GENERIC MAP (
  DEST_SYNC_FF => 2,   -- integer; range: 2-10
  SIM_ASSERT_CHK => 0, -- integer; 0=disable simulation messages, 
                       --          1=enable simulation messages
  SRC_INPUT_REG => 0   -- integer; 0=do not register input, 
                       --          1=register input
)
PORT MAP (
  src_clk => CLK_125MHZ,    -- used only when SRC_INPUT_REG = 1
  src_in => spi_rd_req, 
  dest_clk => CLK_26MHZ,
  dest_out => spi_rd_req_sync
);

-- Acknowledgment of completion of a SPI read request
Sync_spi_rd_ack: xpm_cdc_single
GENERIC MAP (
  DEST_SYNC_FF => 2,   -- integer; range: 2-10
  SIM_ASSERT_CHK => 0, -- integer; 0=disable simulation messages, 
                       --          1=enable simulation messages
  SRC_INPUT_REG => 0   -- integer; 0=do not register input, 
                       --          1=register input
)
PORT MAP (
  src_clk => CLK_26MHZ,    -- used only when SRC_INPUT_REG = 1
  src_in => spi_rd_ack, 
  dest_clk => CLK_125MHZ,
  dest_out => spi_rd_ack_sync
);

--This component is a SERDES (SERializer/DESerializer) circuit
-- that implements a (very) simplified 8-bit SPI (Serial 
-- Peripheral Interface) interface with only two instructions:
-- read and write. See entity comments for further details on
-- operations and I/Os.
SPI_CONTROL_LOGIC: entity work.SPI_MASTER 
PORT MAP(
	CLK => CLK_26MHZ,
	RST => btn_db_26MHZ(0),
	EN_SPI => en_spi_sync,
	PDATA_TO_SPI => pdata_to_spi,
	PDATA_FROM_SPI => pdata_from_spi,
	SPI_SCK => spi_sck_int,
	SPI_S_INV => spi_cs_inv_int,
	SPI_MOSI => spi_mosi_int,
	SPI_MISO => spi_miso_int,
	SPI_WR_REQ => spi_wr_req_sync,
	SPI_WR_ACK => spi_wr_ack,
	SPI_RD_REQ => spi_rd_req_sync,
	SPI_RD_ACK => spi_rd_ack
);

-- Internal signal to I/O mapping (to allow scoping with the ILA)
LED <= LD_INT;
SPI_SCK <= spi_sck_int;
SPI_CS_INV <= spi_cs_inv_int;
SPI_HOLD_INV <= '1';  -- not used in these experiments
SPI_MOSI <= spi_mosi_int;
spi_miso_int <= SPI_MISO; -- not strictly necessary (for completeness only)

-- ChipScope ILA instantiation
-- Note: the first four ports are triggers and might have to be 
--   changed depending on your choice of buttons
-- UNCOMMENT TO USE ILA
ILA: ENTITY work.ila_0
PORT MAP (
  clk => gclk,
  probe0(0) => btn_db_125MHz(0),  -- Reset (BTN0)
  probe1(0) => btn_db_125MHz(1),  -- Pushbutton A (BTN1)
  probe2(0) => btn_db_125MHz(2),  -- Pushbutton B (BTN2)
  probe3(0) => btn_db_125MHz(3),  -- Pushbutton C (BTN3)
  probe4 => LD_INT,
  probe5(0) => spi_sck_int,
  probe6(0) => spi_cs_inv_int,
  probe7(0) => spi_mosi_int,
  probe8(0) => spi_miso_int,
  probe9(0) => spi_hold_inv_int,
  probe10(0) => en_spi,
  probe11(0) => en_spi_sync,
  probe12(0) => spi_wr_req,
  probe13(0) => spi_wr_req_sync,
  probe14(0) => spi_wr_ack,
  probe15(0) => spi_wr_ack_sync,
  probe16 => pdata_to_spi,
  probe17(0) => spi_rd_req,
  probe18(0) => spi_rd_req_sync,
  probe19(0) => spi_rd_ack,
  probe20(0) => spi_rd_ack_sync,
  probe21 => pdata_from_spi
  );

end Behavioral;

